module main

fn main() {
    btree_main()
}
